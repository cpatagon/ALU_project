-- Restador
