-- Divisor
