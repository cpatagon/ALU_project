-- Banco de pruebas del divisor
