-- Paquete de utilidades
