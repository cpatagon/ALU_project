-- Multiplicador
