-- Banco de pruebas del multiplicador
