-- Banco de pruebas del restador
