-- Banco de pruebas del sumador
