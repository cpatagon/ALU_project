-- Multiplexor
